giresh is very good boy
