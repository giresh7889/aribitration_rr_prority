pavan ia doooo
